module tb();
reg clk,rst;
wire Jsel,Jrsel,regwrite,RegDst,ALUsrc,PCSrc,MemRead,MemWrite,MemToReg,zero;
wire [2:0]ALU_operation;
wire [1:0] alu_op;
wire [5:0] OPC,Func;
mips MIPS(clk,rst,Jsel,Jrsel,regwrite,RegDst,ALUsrc,PCSrc,ALU_operation,MemRead,MemWrite,MemToReg,zero,OPC,Func);
controller CONTROLLER(clk,rst,zero,OPC,ALUsrc,Jsel,regwrite,RegDst,alu_op,MemRead,MemWrite,MemToReg,PCSrc);
ALU_controller ALU_CONTROLLER(clk,alu_op,Func,ALU_operation,Jrsel);
initial begin
    #10 rst = 1;
    #20 rst = 0; 
    #20 clk=0;  
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;


end
endmodule